* C:\Users\mayan\eSim-Workspace\AstableMultivibratorUsing555\AstableMultivibratorUsing555.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/07/22 20:15:57

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  GND Capacitor-Voltage OutputVoltage Net-_R1-Pad1_ Net-_C2-Pad1_ Capacitor-Voltage Net-_R1-Pad2_ Net-_R1-Pad1_ LM555N		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 1k		
R2  Net-_R1-Pad2_ Capacitor-Voltage 10k		
C1  Capacitor-Voltage GND 0.1u		
C2  Net-_C2-Pad1_ GND 0.01u		
R3  OutputVoltage GND 1k		
U2  OutputVoltage plot_v1		
U1  Capacitor-Voltage plot_v1		
v1  Net-_R1-Pad1_ GND DC		

.end
